* NGSPICE file created from OR3.ext - technology: scmos

.global Vdd Gnd 

.subckt not gnd VDD in out
M1000 out in gnd Gnd nfet w=2.4u l=1.2u
+  ad=7.2p pd=10.8u as=7.2p ps=10.8u
M1001 out in VDD w_n9_1# pfet w=2.4u l=1.2u
+  ad=7.2p pd=10.8u as=7.2p ps=10.8u
.ends


* Top level circuit OR3

Xnot_0 gnd vdd not_0/in out not
M1000 not_0/in C gnd Gnd nfet w=3.6u l=1.2u
+  ad=66.96p pd=58.8u as=73.44p ps=62.4u
M1001 not_0/in B gnd Gnd nfet w=3.6u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_n42_10# A vdd w_n59_4# pfet w=3.6u l=1.2u
+  ad=54p pd=37.2u as=15.12p ps=15.6u
M1003 not_0/in C a_n15_10# w_n59_4# pfet w=3.6u l=1.2u
+  ad=32.4p pd=25.2u as=66.96p ps=44.4u
M1004 a_n15_10# B a_n42_10# w_n59_4# pfet w=3.6u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
M1005 not_0/in A gnd Gnd nfet w=3.6u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
.end

