magic
tech scmos
timestamp 1701851167
<< metal1 >>
rect 3816 5101 6452 5105
rect 6448 5022 6452 5101
rect 6677 5083 6680 5096
rect 6537 5022 6562 5024
rect 6448 5020 6562 5022
rect 6582 5023 6592 5027
rect 6607 5024 6622 5028
rect 6448 5018 6544 5020
rect 6582 5009 6586 5023
rect 6023 5005 6586 5009
rect 6607 4993 6615 5024
rect 6389 4985 6615 4993
rect 6778 4992 6927 4995
rect 6389 4965 6397 4985
rect 6155 4957 6397 4965
rect 1829 4920 2565 4923
rect 536 4830 1756 4835
rect 536 1881 541 4830
rect 536 1876 1814 1881
rect 536 668 541 1876
rect 1038 1489 1531 1495
rect 1809 1493 1814 1876
rect 811 608 854 611
rect 811 581 814 608
rect 872 604 876 612
rect 1038 605 1044 1489
rect 1829 1449 1832 4920
rect 2562 4843 2565 4920
rect 2562 4840 2693 4843
rect 2743 4825 2805 4830
rect 2833 4825 2845 4830
rect 2743 4806 2748 4825
rect 2698 4801 2748 4806
rect 2633 4758 2655 4762
rect 2563 4757 2655 4758
rect 2563 4753 2638 4757
rect 3746 3736 5764 3740
rect 1734 1446 1832 1449
rect 1890 3519 2383 3522
rect 1504 1439 1522 1444
rect 1586 1443 1593 1445
rect 1580 1442 1593 1443
rect 1580 1440 1589 1442
rect 523 578 814 581
rect 822 600 876 604
rect 983 602 1044 605
rect -88 549 11 553
rect -91 435 9 439
rect 536 406 539 539
rect 822 406 826 600
rect 527 403 826 406
rect 1093 549 1098 1430
rect 526 224 1033 227
rect 507 51 1040 54
rect 387 -240 937 -230
rect 829 -2891 839 -240
rect 829 -2901 959 -2891
rect 1037 -3159 1040 51
rect 1093 -1393 1098 544
rect 1093 -4084 1098 -1398
rect 1093 -4106 1098 -4089
rect 1133 671 1138 1430
rect 1133 -1278 1138 666
rect 1133 -3855 1138 -1283
rect 1133 -4111 1138 -3860
rect 1176 792 1181 1430
rect 1176 -1148 1181 787
rect 1176 -3615 1181 -1153
rect 1176 -4124 1181 -3620
rect 1224 922 1229 1430
rect 1224 -1023 1229 917
rect 1224 -3347 1229 -1028
rect 1224 -4121 1229 -3352
rect 1271 1046 1276 1429
rect 1271 -898 1276 1041
rect 1271 -3996 1276 -903
rect 1271 -4151 1276 -4001
rect 1318 1185 1323 1430
rect 1318 -766 1323 1180
rect 1318 -3743 1323 -771
rect 1318 -4129 1323 -3748
rect 1369 1322 1374 1432
rect 1369 -623 1374 1317
rect 1369 -3478 1374 -628
rect 1369 -4111 1374 -3483
rect 1421 1431 1426 1433
rect 1504 1431 1509 1439
rect 1421 1426 1509 1431
rect 1421 -507 1426 1426
rect 1890 1331 1893 3519
rect 2620 3474 2643 3479
rect 2466 3395 2584 3399
rect 1732 1328 1893 1331
rect 1963 2184 2447 2187
rect 1569 1325 1601 1328
rect 1569 1322 1572 1325
rect 1963 1194 1966 2184
rect 2466 2130 2470 3395
rect 3736 2426 5478 2430
rect 2637 2164 2657 2169
rect 1738 1191 1966 1194
rect 2408 2126 2470 2130
rect 1569 1188 1602 1191
rect 1569 1185 1572 1188
rect 1740 1061 2395 1064
rect 1568 1057 1607 1060
rect 1568 1046 1571 1057
rect 2408 1021 2412 2126
rect 2306 1017 2412 1021
rect 2449 2084 2624 2088
rect 1860 991 1884 995
rect 2209 949 2213 1013
rect 2161 945 2213 949
rect 1571 931 1600 934
rect 1738 933 1894 936
rect 1571 922 1574 931
rect 1891 905 1894 933
rect 1891 902 1938 905
rect 1747 813 1835 816
rect 1566 809 1596 812
rect 1568 792 1571 809
rect 1832 702 1835 813
rect 1865 788 1883 792
rect 2306 746 2310 1017
rect 2449 970 2453 2084
rect 3742 1196 4406 1200
rect 2163 742 2310 746
rect 2348 966 2453 970
rect 2348 704 2352 966
rect 2554 940 2561 1062
rect 2554 933 2691 940
rect 3959 900 4042 903
rect 1832 699 1937 702
rect 2214 700 2352 704
rect 2426 852 2653 856
rect 1751 682 1835 685
rect 1566 678 1595 681
rect 1568 671 1571 678
rect 1762 562 1779 565
rect 1572 559 1594 562
rect 1568 556 1575 559
rect 1776 172 1779 562
rect 1832 464 1835 682
rect 1858 549 1881 553
rect 2214 507 2218 700
rect 2160 503 2218 507
rect 1832 461 1932 464
rect 1854 273 1883 277
rect 1854 262 1858 273
rect 1830 258 1858 262
rect 1879 259 1883 273
rect 2426 217 2430 852
rect 2163 213 2430 217
rect 1776 169 1937 172
rect 2784 21 2868 31
rect 2784 -67 2794 21
rect 1861 -77 2794 -67
rect 1861 -230 1871 -77
rect 4402 -145 4406 1196
rect 5474 -29 5478 2426
rect 5760 992 5764 3736
rect 5760 988 6048 992
rect 5474 -33 6073 -29
rect 4402 -149 6122 -145
rect 1465 -240 1871 -230
rect 2020 -154 2337 -151
rect 1785 -269 1793 -240
rect 1537 -462 1576 -457
rect 2020 -502 2023 -154
rect 2334 -161 2337 -154
rect 2364 -161 2402 -159
rect 2334 -162 2402 -161
rect 2334 -164 2367 -162
rect 5001 -237 5224 -231
rect 2403 -243 2429 -240
rect 2403 -246 2406 -243
rect 2426 -252 2429 -243
rect 5218 -278 5224 -237
rect 5129 -286 5156 -283
rect 5153 -339 5156 -286
rect 5557 -314 5593 -311
rect 5153 -342 5184 -339
rect 5199 -348 5202 -339
rect 5557 -343 5560 -314
rect 5291 -346 5560 -343
rect 5156 -351 5202 -348
rect 4040 -472 6092 -469
rect 1781 -505 2023 -502
rect 1421 -512 1575 -507
rect 1634 -508 1640 -506
rect 1626 -509 1640 -508
rect 1626 -511 1637 -509
rect 1421 -3222 1426 -512
rect 2332 -587 2365 -584
rect 2332 -620 2335 -587
rect 1779 -623 2335 -620
rect 1612 -626 1650 -623
rect 5210 -657 5215 -531
rect 4981 -662 5215 -657
rect 4981 -663 4986 -662
rect 2427 -676 2448 -673
rect 2235 -685 2362 -680
rect 1786 -760 2324 -757
rect 1607 -763 1649 -760
rect 1607 -766 1610 -763
rect 1787 -890 2230 -887
rect 1606 -894 1654 -891
rect 1606 -898 1609 -894
rect 2043 -1015 2046 -917
rect 1607 -1020 1649 -1017
rect 1785 -1018 2046 -1015
rect 2118 -934 2165 -931
rect 1607 -1023 1610 -1020
rect 2118 -1135 2121 -934
rect 1795 -1138 2121 -1135
rect 2179 -1133 2193 -1130
rect 1609 -1142 1644 -1139
rect 1609 -1148 1612 -1142
rect 2179 -1266 2182 -1133
rect 1797 -1269 2182 -1266
rect 1610 -1273 1641 -1270
rect 1610 -1278 1613 -1273
rect 1810 -1389 2146 -1386
rect 1553 -1392 1641 -1389
rect 1553 -1393 1556 -1392
rect 1537 -1396 1556 -1393
rect 2143 -1588 2146 -1389
rect 2227 -1504 2230 -890
rect 2321 -1041 2324 -760
rect 3701 -827 3704 -818
rect 3918 -825 3952 -822
rect 3957 -825 4305 -820
rect 5865 -825 6116 -820
rect 3705 -839 3708 -832
rect 2321 -1044 2358 -1041
rect 2321 -1046 2324 -1044
rect 2256 -1134 2312 -1129
rect 2419 -1134 2436 -1131
rect 4126 -1367 4278 -1364
rect 2227 -1507 2312 -1504
rect 6155 -1540 6163 4957
rect 6647 4915 6652 4938
rect 6591 4910 6652 4915
rect 6591 3978 6596 4910
rect 6591 3973 9022 3978
rect 7507 887 7512 914
rect 7204 883 7266 887
rect 7176 833 7193 837
rect 7189 816 7193 833
rect 7262 832 7266 883
rect 7262 828 7430 832
rect 7450 831 7460 835
rect 7481 832 7490 836
rect 7450 816 7454 831
rect 7189 812 7454 816
rect 7481 796 7484 832
rect 7649 800 7809 803
rect 7347 793 7484 796
rect 7347 754 7350 793
rect 6888 751 7350 754
rect 6711 -33 6823 -26
rect 6690 -149 6823 -143
rect 6719 -472 6862 -466
rect 5476 -1543 6163 -1540
rect 2143 -1591 2299 -1588
rect 2401 -1589 2415 -1586
rect 2412 -1595 2415 -1589
rect 1571 -3180 1633 -3175
rect 1838 -3222 2230 -3219
rect 1678 -3226 1697 -3223
rect 1421 -4116 1426 -3227
rect 2227 -3249 2230 -3222
rect 2227 -3252 2265 -3249
rect 2280 -3257 2283 -3249
rect 5476 -3253 5479 -1543
rect 6155 -1545 6163 -1543
rect 2372 -3256 5479 -3253
rect 1935 -3260 2283 -3257
rect 1935 -3337 1938 -3260
rect 1836 -3340 1938 -3337
rect 1671 -3343 1705 -3340
rect 1671 -3347 1674 -3343
rect 1844 -3477 2245 -3474
rect 1673 -3488 1676 -3483
rect 1703 -3488 1706 -3477
rect 1673 -3491 1706 -3488
rect 2242 -3499 2245 -3477
rect 2242 -3502 2270 -3499
rect 2285 -3505 2288 -3499
rect 6888 -3503 6891 751
rect 7503 14 7508 745
rect 9017 14 9022 3973
rect 7503 9 10425 14
rect 9521 -632 9560 -628
rect 9556 -662 9560 -632
rect 9556 -666 9774 -662
rect 10032 -666 10035 -636
rect 9770 -725 9774 -666
rect 9770 -729 9886 -725
rect 9907 -726 9916 -722
rect 9934 -725 9946 -721
rect 9611 -737 9627 -733
rect 9623 -746 9627 -737
rect 9907 -746 9911 -726
rect 9623 -750 9911 -746
rect 9934 -761 9938 -725
rect 10105 -757 10278 -754
rect 9691 -765 9938 -761
rect 9691 -799 9695 -765
rect 9666 -800 9695 -799
rect 1937 -3508 2288 -3505
rect 2377 -3506 6891 -3503
rect 8452 -803 9695 -800
rect 1937 -3604 1940 -3508
rect 1838 -3607 1940 -3604
rect 1671 -3611 1711 -3608
rect 1671 -3615 1674 -3611
rect 2222 -3722 2266 -3719
rect 2222 -3732 2225 -3722
rect 2282 -3726 2285 -3719
rect 8452 -3723 8455 -803
rect 9978 -863 9983 -811
rect 10420 -863 10425 9
rect 9978 -868 10425 -863
rect 9978 -989 9983 -868
rect 9756 -994 9983 -989
rect 9756 -2040 9761 -994
rect 10795 -1913 10845 -1909
rect 10841 -2003 10845 -1913
rect 10841 -2007 11364 -2003
rect 11382 -2012 11385 -2003
rect 11346 -2015 11385 -2012
rect 11493 -2013 11587 -2010
rect 11346 -2028 11349 -2015
rect 11177 -2031 11349 -2028
rect 11177 -2055 11180 -2031
rect 2373 -3726 8455 -3723
rect 10140 -2058 11180 -2055
rect 1667 -3737 1704 -3734
rect 1842 -3735 2225 -3732
rect 2244 -3729 2285 -3726
rect 1667 -3743 1670 -3737
rect 2244 -3844 2247 -3729
rect 1864 -3847 2247 -3844
rect 1864 -3852 1867 -3847
rect 1851 -3855 1867 -3852
rect 1675 -3859 1701 -3856
rect 1855 -3985 2234 -3983
rect 1855 -3986 2268 -3985
rect 1671 -3990 1698 -3987
rect 2231 -3988 2268 -3986
rect 1671 -3996 1674 -3990
rect 2284 -3992 2287 -3985
rect 10140 -3989 10143 -2058
rect 2376 -3992 10143 -3989
rect 2055 -3995 2287 -3992
rect 2055 -4103 2058 -3995
rect 1863 -4106 2058 -4103
rect 1626 -4115 1629 -4113
rect 1646 -4109 1698 -4106
rect 1646 -4115 1649 -4109
rect 1626 -4118 1649 -4115
<< m2contact >>
rect 6677 5096 6682 5101
rect 6018 5005 6023 5010
rect 1756 4830 1761 4835
rect 536 663 541 668
rect 1809 1488 1814 1493
rect 2805 4825 2810 4830
rect 2828 4825 2833 4830
rect 2693 4801 2698 4806
rect 2558 4753 2563 4758
rect 1522 1439 1527 1444
rect 1575 1439 1580 1444
rect 536 539 541 544
rect 1093 544 1098 549
rect 1033 224 1038 229
rect 377 -240 387 -230
rect 937 -240 947 -230
rect 959 -2901 974 -2886
rect 1093 -1398 1098 -1393
rect 1037 -3164 1043 -3159
rect 1093 -4089 1098 -4084
rect 1133 666 1138 671
rect 1133 -1283 1138 -1278
rect 1133 -3860 1138 -3855
rect 1176 787 1181 792
rect 1176 -1153 1181 -1148
rect 1176 -3620 1181 -3615
rect 1224 917 1229 922
rect 1224 -1028 1229 -1023
rect 1224 -3352 1229 -3347
rect 1271 1041 1276 1046
rect 1271 -903 1276 -898
rect 1271 -4001 1276 -3996
rect 1318 1180 1323 1185
rect 1318 -771 1323 -766
rect 1318 -3748 1323 -3743
rect 1369 1317 1374 1322
rect 1369 -628 1374 -623
rect 1369 -3483 1374 -3478
rect 2383 3517 2388 3522
rect 2615 3474 2620 3479
rect 1567 1317 1572 1322
rect 2447 2182 2452 2187
rect 2632 2164 2637 2169
rect 1568 1180 1573 1185
rect 2395 1058 2401 1064
rect 1567 1041 1572 1046
rect 2209 1013 2214 1018
rect 1855 990 1860 995
rect 1570 917 1575 922
rect 1567 787 1572 792
rect 1860 787 1865 792
rect 2554 1062 2561 1069
rect 1567 666 1572 671
rect 1563 556 1568 561
rect 1853 549 1858 554
rect 1825 257 1830 262
rect 2868 21 2878 31
rect 6048 988 6055 995
rect 6073 -33 6080 -26
rect 6122 -149 6128 -143
rect 1455 -240 1465 -230
rect 1785 -278 1793 -269
rect 1532 -462 1537 -457
rect 4995 -237 5001 -231
rect 2403 -251 2408 -246
rect 5124 -286 5129 -281
rect 5218 -284 5224 -278
rect 5593 -315 5598 -310
rect 5151 -353 5156 -348
rect 6092 -472 6098 -466
rect 1575 -512 1580 -507
rect 1621 -512 1626 -507
rect 5210 -531 5215 -526
rect 1607 -628 1612 -623
rect 4976 -663 4981 -657
rect 2422 -678 2427 -673
rect 2230 -685 2235 -680
rect 2362 -685 2367 -680
rect 1606 -771 1611 -766
rect 1605 -903 1610 -898
rect 2043 -917 2048 -912
rect 2165 -934 2170 -929
rect 1607 -1028 1612 -1023
rect 1607 -1153 1612 -1148
rect 2193 -1134 2198 -1129
rect 1609 -1283 1614 -1278
rect 1532 -1398 1537 -1393
rect 3952 -825 3957 -820
rect 4305 -825 4310 -820
rect 5860 -825 5865 -820
rect 6116 -825 6121 -820
rect 2251 -1134 2256 -1129
rect 2312 -1134 2317 -1129
rect 2414 -1134 2419 -1129
rect 4278 -1367 4283 -1362
rect 7507 914 7512 919
rect 7197 881 7204 888
rect 7171 833 7176 838
rect 6704 -33 6711 -26
rect 6823 -33 6830 -26
rect 6684 -149 6690 -143
rect 6823 -149 6829 -143
rect 6713 -472 6719 -466
rect 6862 -472 6868 -466
rect 2299 -1591 2304 -1586
rect 2396 -1591 2401 -1586
rect 1566 -3180 1571 -3175
rect 1421 -3227 1426 -3222
rect 1673 -3227 1678 -3222
rect 1670 -3352 1675 -3347
rect 1672 -3483 1677 -3478
rect 9514 -633 9521 -626
rect 10031 -636 10036 -631
rect 9605 -737 9611 -731
rect 1670 -3620 1675 -3615
rect 10789 -1915 10795 -1909
rect 9756 -2045 9761 -2040
rect 1666 -3748 1671 -3743
rect 1670 -3860 1675 -3855
rect 1670 -4001 1675 -3996
rect 1624 -4113 1629 -4108
<< metal2 >>
rect 474 5972 3458 5973
rect 474 5968 6682 5972
rect 474 1793 479 5968
rect 3453 5967 6682 5968
rect 3453 5330 3458 5967
rect 6677 5101 6682 5967
rect 6682 5096 6879 5101
rect 5959 5005 6018 5010
rect 1761 4830 2538 4835
rect 2533 4806 2538 4830
rect 2810 4825 2828 4830
rect 2533 4801 2693 4806
rect 2209 4753 2558 4758
rect 474 1788 1727 1793
rect 474 701 479 1788
rect 1722 1539 1727 1788
rect 1783 1530 1998 1535
rect 1527 1439 1575 1444
rect 1374 1317 1567 1322
rect 1323 1180 1568 1185
rect 1276 1041 1567 1046
rect 1809 995 1814 1488
rect 1993 1091 1998 1530
rect 1878 1086 1998 1091
rect 1809 990 1855 995
rect 1229 917 1570 922
rect 1809 792 1814 990
rect 1878 852 1883 1086
rect 1993 1031 1998 1086
rect 2209 1018 2214 4753
rect 2388 3517 2620 3522
rect 2615 3479 2620 3517
rect 2452 2182 2637 2187
rect 2632 2169 2637 2182
rect 2537 1072 2560 1078
rect 2537 1064 2543 1072
rect 2401 1058 2543 1064
rect 2554 1069 2560 1072
rect 2099 864 2107 882
rect 2099 856 2199 864
rect 1878 847 2019 852
rect 1181 787 1567 792
rect 1809 787 1860 792
rect 474 696 860 701
rect -11 663 117 668
rect 474 663 479 696
rect -11 -235 -6 663
rect 536 544 541 663
rect 855 656 860 696
rect 1138 666 1567 671
rect 916 469 924 558
rect 1563 549 1568 556
rect 1098 544 1568 549
rect 1809 554 1814 787
rect 1878 626 1883 847
rect 2014 828 2019 847
rect 2096 663 2104 677
rect 2191 663 2199 856
rect 2096 655 2199 663
rect 1878 621 2008 626
rect 1809 549 1853 554
rect 589 464 924 469
rect 589 5 594 464
rect 916 441 924 464
rect 1609 462 1617 511
rect 1609 454 1690 462
rect 1642 441 1650 454
rect 916 433 1650 441
rect 1038 224 1537 229
rect 338 0 594 5
rect -11 -240 377 -235
rect 506 -2522 511 0
rect 1532 -55 1537 224
rect 1682 -2 1690 454
rect 1809 262 1814 549
rect 1878 357 1883 621
rect 2003 590 2008 621
rect 2089 404 2097 439
rect 2191 404 2199 655
rect 2247 495 2291 503
rect 2089 396 2201 404
rect 1878 352 2012 357
rect 2007 299 2012 352
rect 1809 257 1825 262
rect 2079 81 2087 150
rect 2193 81 2201 396
rect 2079 73 2201 81
rect 2079 -2 2087 73
rect 2502 -2 2510 502
rect 1682 -10 2510 -2
rect 2668 237 5062 242
rect 2668 -43 2673 237
rect 1819 -48 2673 -43
rect 1819 -55 1824 -48
rect 1532 -60 1824 -55
rect 947 -240 1455 -230
rect 1532 -457 1537 -60
rect 2872 -66 2876 21
rect 4889 -237 4995 -231
rect 2403 -259 2408 -251
rect 2188 -264 2408 -259
rect 1785 -413 1790 -278
rect 1580 -512 1621 -507
rect 2188 -570 2193 -264
rect 4889 -345 4895 -237
rect 5057 -281 5062 237
rect 5057 -286 5124 -281
rect 5598 -315 5728 -310
rect 4092 -351 4895 -345
rect 2043 -575 2193 -570
rect 5052 -353 5151 -348
rect 1374 -628 1607 -623
rect 1323 -771 1606 -766
rect 1276 -903 1605 -898
rect 2043 -912 2048 -575
rect 4208 -663 4976 -660
rect 2422 -680 2427 -678
rect 2165 -685 2230 -680
rect 2367 -685 2427 -680
rect 2165 -929 2170 -685
rect 5052 -820 5057 -353
rect 5215 -505 5220 -364
rect 5209 -510 5220 -505
rect 5209 -526 5214 -510
rect 5209 -528 5210 -526
rect 5723 -820 5728 -315
rect 4310 -825 5058 -820
rect 5722 -825 5860 -820
rect 3769 -866 3781 -862
rect 3789 -870 3801 -867
rect 1229 -1028 1607 -1023
rect 2198 -1134 2251 -1129
rect 2317 -1134 2414 -1129
rect 1181 -1153 1607 -1148
rect 1630 -1200 1635 -1159
rect 1138 -1283 1609 -1278
rect 5959 -1362 5964 5005
rect 6874 1138 6879 5096
rect 6874 1133 7697 1138
rect 6055 988 6649 995
rect 6642 888 6649 988
rect 7507 919 7512 1133
rect 6642 881 7197 888
rect 6755 833 7171 838
rect 6080 -33 6704 -26
rect 6128 -149 6684 -143
rect 6098 -472 6713 -466
rect 6755 -820 6760 833
rect 7692 312 7697 1133
rect 7692 307 10152 312
rect 6830 -33 8577 -26
rect 6121 -825 6760 -820
rect 6829 -979 6835 -143
rect 6868 -472 8081 -466
rect 8075 -731 8081 -472
rect 8570 -626 8577 -33
rect 10147 -599 10152 307
rect 10031 -604 10152 -599
rect 8570 -633 9514 -626
rect 10031 -631 10036 -604
rect 8075 -737 9605 -731
rect 6829 -985 7086 -979
rect 4283 -1367 5964 -1362
rect 1098 -1398 1532 -1393
rect 1674 -1709 1678 -1437
rect 2304 -1591 2396 -1586
rect 1674 -1713 2270 -1709
rect 7080 -2014 7086 -985
rect 10147 -1496 10152 -604
rect 10147 -1501 11403 -1496
rect 9949 -1915 10789 -1909
rect 9949 -2014 9955 -1915
rect 11398 -1957 11403 -1501
rect 7080 -2020 9955 -2014
rect 2438 -2522 2443 -2068
rect 9756 -2139 9761 -2045
rect 11432 -2139 11437 -2061
rect 9756 -2144 11437 -2139
rect 506 -2527 2443 -2522
rect 735 -4200 740 -2527
rect 974 -2901 1843 -2886
rect 1828 -3078 1843 -2901
rect 1828 -3093 2180 -3078
rect 1828 -3127 1843 -3093
rect 2165 -3152 2180 -3093
rect 2165 -3157 2293 -3152
rect 1043 -3164 1571 -3159
rect 1566 -3175 1571 -3164
rect 1426 -3227 1673 -3222
rect 1229 -3352 1670 -3347
rect 2165 -3409 2180 -3157
rect 2288 -3199 2293 -3157
rect 2309 -3329 2314 -3277
rect 2309 -3334 2429 -3329
rect 2165 -3414 2309 -3409
rect 1374 -3483 1672 -3478
rect 1181 -3620 1670 -3615
rect 2165 -3631 2180 -3414
rect 2304 -3449 2309 -3414
rect 2312 -3568 2317 -3524
rect 2424 -3568 2429 -3334
rect 2312 -3573 2429 -3568
rect 2165 -3636 2304 -3631
rect 1323 -3748 1666 -3743
rect 1138 -3860 1670 -3855
rect 2165 -3911 2180 -3636
rect 2299 -3669 2304 -3636
rect 2311 -3834 2316 -3744
rect 2424 -3834 2429 -3573
rect 2311 -3839 2429 -3834
rect 2165 -3916 2295 -3911
rect 2165 -3920 2180 -3916
rect 2290 -3935 2295 -3916
rect 1276 -4001 1670 -3996
rect 1098 -4089 1629 -4084
rect 1624 -4108 1629 -4089
rect 2320 -4152 2325 -4013
rect 2424 -4152 2429 -3839
rect 2320 -4155 2429 -4152
rect 1507 -4161 1696 -4156
rect 1730 -4157 2429 -4155
rect 1730 -4160 2325 -4157
rect 1507 -4198 1512 -4161
rect 11432 -4198 11437 -2144
rect 1507 -4200 11437 -4198
rect 735 -4203 11437 -4200
rect 735 -4205 1512 -4203
use OR  OR_0
timestamp 1701543975
transform 1 0 854 0 1 571
box -4 -21 132 92
use XOR  XOR_3
timestamp 1701356350
transform 1 0 2015 0 1 235
box -136 -88 152 66
use XOR  XOR_2
timestamp 1701356350
transform 1 0 2012 0 1 525
box -136 -88 152 66
use decoder  decoder_0
timestamp 1701836177
transform 1 0 108 0 1 534
box -108 -534 423 134
use enable  enable_0
timestamp 1701538289
transform 1 0 1613 0 1 1423
box -89 -916 175 120
use enable  enable_1
timestamp 1701538289
transform 1 0 1660 0 1 -528
box -89 -916 175 120
use enable  enable_2
timestamp 1701538289
transform 1 0 1717 0 1 -3245
box -89 -916 175 120
use XOR  XOR_0
timestamp 1701356350
transform 1 0 2014 0 1 967
box -136 -88 152 66
use XOR  XOR_1
timestamp 1701356350
transform 1 0 2015 0 1 764
box -136 -88 152 66
use four_bit_adder  four_bit_adder_0
timestamp 1701849322
transform 1 0 2673 0 1 4636
box -406 -4141 1643 698
use AND  AND_3
timestamp 1701359634
transform 1 0 2268 0 1 -4011
box -2 -4 111 81
use AND  AND_2
timestamp 1701359634
transform 1 0 2266 0 1 -3745
box -2 -4 111 81
use AND  AND_1
timestamp 1701359634
transform 1 0 2269 0 1 -3525
box -2 -4 111 81
use AND  AND_0
timestamp 1701359634
transform 1 0 2264 0 1 -3275
box -2 -4 111 81
use comparator  comparator_0
timestamp 1701502639
transform 1 0 2509 0 1 -293
box -243 -1779 1831 231
use AND  AND_4
timestamp 1701359634
transform 1 0 5183 0 1 -365
box -2 -4 111 81
use OR3  OR3_1
timestamp 1701521602
transform 1 0 7485 0 1 863
box -59 -123 167 31
use OR3  OR3_0
timestamp 1701521602
transform 1 0 6617 0 1 5055
box -59 -123 167 31
use OR3  OR3_2
timestamp 1701521602
transform 1 0 9941 0 1 -694
box -59 -123 167 31
use OR  OR_1
timestamp 1701543975
transform 1 0 11364 0 1 -2044
box -4 -21 132 92
<< labels >>
rlabel metal1 -85 436 -83 437 1 S1
rlabel metal1 -77 550 -75 551 1 S0
rlabel metal1 556 579 558 580 1 en0
rlabel metal1 573 404 575 405 1 en1
rlabel metal1 570 225 572 226 1 en2
rlabel metal1 573 52 575 53 1 en3
rlabel metal1 1423 1427 1425 1429 1 A0
rlabel metal1 1371 1428 1373 1430 1 A1
rlabel metal1 1319 1425 1321 1427 1 A2
rlabel metal1 1272 1424 1274 1426 1 A3
rlabel metal1 1225 1425 1227 1427 1 B0
rlabel metal1 1177 1425 1179 1427 1 B1
rlabel metal1 1135 1425 1137 1427 1 B2
rlabel metal1 1095 1425 1097 1427 1 B3
rlabel metal1 6924 4993 6926 4994 1 Out0
rlabel metal1 7795 801 7797 802 1 Out1
rlabel metal1 10271 -756 10273 -755 1 Out2
rlabel metal1 11580 -2012 11583 -2011 1 Out3
rlabel metal1 4035 901 4038 902 1 Out4
rlabel metal2 1241 -4204 1245 -4203 1 gnd
rlabel metal2 3701 5969 3708 5970 5 vdd
rlabel metal2 7080 883 7084 885 1 outout1
rlabel metal2 7081 834 7085 836 1 outout2
rlabel metal1 7100 752 7104 754 1 outout3
rlabel metal1 3933 -824 3936 -823 1 eequal
rlabel space 3695 -826 3698 -825 1 ea1
rlabel space 3760 -882 3763 -881 1 ea3
rlabel space 3697 -834 3700 -833 1 ea2
rlabel space 3774 -922 3777 -921 1 ea4
rlabel metal1 3702 -821 3703 -820 1 ea1
rlabel metal1 3706 -838 3707 -837 1 ea2
rlabel metal2 3770 -865 3771 -864 1 ea3
rlabel metal2 3790 -869 3792 -868 1 ea4
rlabel metal1 1898 -504 1900 -503 1 f0
rlabel metal1 1915 -623 1917 -622 1 f1
rlabel metal1 1913 -759 1915 -758 1 f2
rlabel metal1 1912 -889 1914 -888 1 f3
rlabel metal1 1915 -1018 1917 -1017 1 f4
rlabel metal1 1912 -1137 1914 -1136 1 f5
rlabel metal1 1919 -1268 1921 -1267 1 f6
rlabel metal1 1935 -1388 1937 -1387 1 f7
<< end >>
