* NGSPICE file created from AND4.ext - technology: scmos

.global Vdd Gnd 

.subckt not gnd VDD in out
M1000 out in gnd Gnd nfet w=2.4u l=1.2u
+  ad=7.2p pd=10.8u as=7.2p ps=10.8u
M1001 out in VDD w_n9_1# pfet w=2.4u l=1.2u
+  ad=7.2p pd=10.8u as=7.2p ps=10.8u
.ends


* Top level circuit AND4

Xnot_0 gnd vdd not_0/in out not
M1000 not_0/in D a_25_n36# Gnd nfet w=3u l=1.2u
+  ad=14.4p pd=15.6u as=30.6p ps=26.4u
M1001 a_6_n36# B a_n14_n36# Gnd nfet w=3u l=1.2u
+  ad=30.6p pd=26.4u as=32.4p ps=27.6u
M1002 not_0/in D vdd w_n27_2# pfet w=3u l=1.2u
+  ad=37.8p pd=49.2u as=41.4p ps=51.6u
M1003 not_0/in C vdd w_n27_2# pfet w=3u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_25_n36# C a_6_n36# Gnd nfet w=3u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_n14_n36# A gnd Gnd nfet w=3u l=1.2u
+  ad=0p pd=0u as=14.4p ps=15.6u
M1006 not_0/in B vdd w_n27_2# pfet w=3u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
M1007 not_0/in A vdd w_n27_2# pfet w=3u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
.end

