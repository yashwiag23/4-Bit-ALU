magic
tech scmos
timestamp 1701502639
<< metal1 >>
rect -122 130 6 134
rect -95 101 -91 130
rect -140 97 -91 101
rect -140 -99 -136 97
rect 453 87 1045 90
rect -83 41 41 44
rect -48 -43 -45 41
rect 113 -12 626 -6
rect 113 -25 119 -12
rect 153 -22 159 -12
rect 620 -29 626 -12
rect 648 -28 652 -5
rect 756 -34 970 -31
rect -48 -46 144 -43
rect 164 -46 560 -43
rect -4 -63 -1 -46
rect 156 -76 159 -58
rect 156 -79 440 -76
rect 557 -83 560 -46
rect 557 -86 592 -83
rect 606 -91 610 -82
rect 536 -95 610 -91
rect 536 -99 540 -95
rect -140 -103 540 -99
rect -140 -140 -136 -103
rect 119 -118 161 -115
rect 158 -125 161 -118
rect -140 -143 119 -140
rect -140 -144 147 -143
rect 218 -144 586 -140
rect 115 -145 147 -144
rect 115 -148 145 -145
rect 166 -147 222 -144
rect 201 -148 222 -147
rect 115 -151 119 -148
rect 51 -221 57 -170
rect 221 -185 493 -182
rect 490 -258 493 -185
rect 582 -242 586 -144
rect 802 -158 806 -105
rect 855 -194 938 -191
rect 582 -246 693 -242
rect 705 -251 708 -242
rect 661 -254 708 -251
rect 661 -258 664 -254
rect 490 -261 664 -258
rect -157 -294 -5 -290
rect -74 -328 -70 -294
rect -125 -332 -70 -328
rect -125 -516 -121 -332
rect 624 -334 627 -304
rect 699 -318 704 -276
rect 724 -334 727 -286
rect 445 -337 896 -334
rect -64 -383 32 -380
rect -39 -486 -36 -383
rect 828 -466 880 -463
rect -39 -489 145 -486
rect 166 -489 470 -486
rect 13 -496 16 -489
rect 467 -496 470 -489
rect 828 -493 831 -466
rect 630 -496 831 -493
rect 467 -499 479 -496
rect 494 -505 498 -496
rect 435 -509 498 -505
rect 435 -516 439 -509
rect -125 -520 439 -516
rect -125 -589 -121 -520
rect 486 -546 489 -528
rect 893 -539 896 -337
rect 906 -466 995 -463
rect 1042 -515 1045 87
rect 1262 -177 1285 -174
rect 1262 -294 1265 -177
rect 1456 -179 1534 -176
rect 1363 -235 1366 -214
rect 1554 -231 1641 -228
rect 1554 -235 1557 -231
rect 1363 -238 1557 -235
rect 1262 -297 1831 -294
rect 1301 -469 1547 -463
rect 1301 -486 1307 -469
rect 1042 -518 1121 -515
rect 1118 -531 1121 -518
rect 1118 -534 1231 -531
rect 1383 -532 1413 -529
rect 1252 -539 1255 -535
rect 893 -542 1255 -539
rect 294 -549 489 -546
rect 1268 -544 1272 -532
rect 1284 -536 1291 -532
rect 1284 -540 1288 -536
rect 1284 -544 1294 -540
rect 501 -565 628 -560
rect 623 -583 628 -565
rect 1340 -573 1345 -563
rect 1372 -572 1653 -567
rect 1372 -573 1377 -572
rect 1340 -578 1377 -573
rect 130 -589 147 -588
rect -125 -590 147 -589
rect -125 -593 146 -590
rect 166 -592 579 -589
rect 109 -624 112 -609
rect 145 -624 148 -604
rect 109 -627 148 -624
rect 576 -623 579 -592
rect 1206 -621 1209 -612
rect 576 -626 622 -623
rect 145 -652 148 -627
rect 637 -635 640 -624
rect 769 -624 1209 -621
rect 1289 -627 1292 -585
rect 590 -638 640 -635
rect 1239 -630 1292 -627
rect 590 -645 593 -638
rect 463 -648 593 -645
rect 145 -655 150 -652
rect 147 -662 150 -655
rect 623 -664 627 -656
rect 152 -668 627 -664
rect 1239 -666 1242 -630
rect 927 -669 1242 -666
rect 1239 -694 1242 -669
rect 1075 -697 1242 -694
rect -162 -752 -14 -748
rect -111 -1043 -107 -752
rect 431 -795 724 -792
rect -76 -841 24 -838
rect -43 -939 -40 -841
rect 676 -897 773 -891
rect 543 -901 565 -898
rect 543 -914 546 -901
rect 562 -910 565 -901
rect 152 -917 546 -914
rect 676 -915 682 -897
rect 152 -928 155 -917
rect 767 -918 773 -897
rect -43 -942 120 -939
rect 40 -960 43 -942
rect 117 -946 120 -942
rect 117 -949 140 -946
rect 537 -947 558 -945
rect 160 -948 558 -947
rect 160 -950 540 -948
rect 573 -949 580 -945
rect 710 -947 1178 -944
rect 573 -956 577 -949
rect 523 -960 577 -956
rect 523 -994 527 -960
rect 6 -998 527 -994
rect 6 -1043 10 -998
rect 771 -1011 777 -1002
rect 143 -1017 777 -1011
rect 143 -1023 149 -1017
rect 771 -1042 777 -1017
rect -111 -1047 141 -1043
rect 162 -1047 655 -1044
rect 84 -1073 88 -1064
rect 142 -1073 146 -1062
rect 652 -1073 655 -1047
rect 84 -1077 528 -1073
rect 652 -1076 728 -1073
rect 524 -1142 528 -1077
rect 743 -1077 750 -1072
rect 883 -1074 1195 -1071
rect 743 -1083 746 -1077
rect 639 -1086 746 -1083
rect 639 -1091 642 -1086
rect 545 -1094 642 -1091
rect 735 -1142 739 -1107
rect 524 -1146 739 -1142
rect -206 -1213 -6 -1209
rect -173 -1563 -169 -1213
rect -145 -1478 -141 -1213
rect 553 -1240 556 -1146
rect 615 -1253 618 -1190
rect 1239 -1253 1242 -697
rect 1297 -1059 1300 -909
rect 1345 -1053 1348 -910
rect 1345 -1056 1477 -1053
rect 1297 -1062 1455 -1059
rect 1397 -1072 1419 -1069
rect 1433 -1078 1436 -1069
rect 1452 -1075 1455 -1062
rect 1474 -1074 1477 -1056
rect 1590 -1074 1621 -1071
rect 1390 -1081 1436 -1078
rect 1390 -1142 1393 -1081
rect 439 -1256 1242 -1253
rect -97 -1302 26 -1299
rect -73 -1441 -70 -1302
rect -35 -1351 -32 -1302
rect 183 -1441 222 -1440
rect -73 -1444 121 -1441
rect 140 -1443 222 -1441
rect 140 -1444 187 -1443
rect 219 -1474 222 -1443
rect 219 -1477 238 -1474
rect -145 -1481 213 -1478
rect 253 -1481 257 -1475
rect 1828 -1478 1831 -297
rect 345 -1481 1831 -1478
rect -145 -1482 257 -1481
rect 209 -1485 257 -1482
rect -173 -1567 122 -1563
rect 142 -1566 194 -1563
rect 191 -1592 194 -1566
rect 191 -1595 241 -1592
rect 258 -1600 261 -1592
rect 1390 -1596 1393 -1528
rect 350 -1599 1393 -1596
rect 173 -1603 261 -1600
rect 173 -1611 176 -1603
rect -14 -1614 176 -1611
<< m2contact >>
rect 648 -5 654 1
rect 113 -31 119 -25
rect 970 -36 975 -31
rect -4 -68 1 -63
rect 440 -81 445 -76
rect 624 -85 629 -80
rect 644 -86 649 -81
rect 663 -86 668 -81
rect 801 -105 806 -100
rect 113 -118 119 -112
rect 600 -123 606 -117
rect 51 -170 57 -164
rect 158 -167 163 -162
rect 216 -185 221 -180
rect 51 -228 58 -221
rect 938 -194 943 -189
rect 722 -246 727 -241
rect 742 -246 747 -241
rect 761 -247 766 -242
rect 622 -304 627 -299
rect 722 -286 727 -281
rect 699 -323 704 -318
rect 539 -449 544 -444
rect 150 -464 155 -459
rect 880 -466 885 -461
rect 13 -501 18 -496
rect 146 -509 151 -504
rect 511 -501 516 -496
rect 530 -501 535 -496
rect 289 -549 294 -544
rect 901 -466 906 -461
rect 995 -466 1000 -461
rect 1391 -117 1396 -112
rect 1298 -179 1303 -174
rect 1317 -180 1322 -175
rect 1338 -180 1343 -175
rect 1641 -232 1646 -227
rect 1547 -474 1559 -462
rect 1268 -549 1273 -544
rect 1289 -549 1294 -544
rect 146 -567 151 -562
rect 493 -565 501 -557
rect 1653 -572 1665 -560
rect 1289 -585 1294 -580
rect 109 -609 114 -604
rect 1206 -612 1211 -607
rect 653 -629 658 -624
rect 672 -628 677 -623
rect 458 -648 463 -643
rect 146 -668 152 -662
rect 922 -669 927 -664
rect 1070 -697 1075 -692
rect 724 -796 729 -791
rect 476 -914 482 -908
rect 767 -924 773 -918
rect 593 -949 598 -944
rect 1178 -947 1183 -942
rect 40 -965 45 -960
rect 141 -970 147 -965
rect 559 -990 565 -984
rect 771 -1002 777 -996
rect 84 -1064 90 -1058
rect 763 -1077 768 -1072
rect 1195 -1074 1200 -1069
rect 540 -1094 545 -1089
rect 615 -1190 620 -1185
rect 553 -1245 558 -1240
rect 1297 -909 1302 -904
rect 1345 -910 1350 -905
rect 1493 -1012 1502 -1003
rect 1392 -1074 1397 -1069
rect 1508 -1117 1513 -1112
rect 1390 -1147 1395 -1142
rect -35 -1356 -30 -1351
rect 119 -1419 124 -1414
rect 119 -1464 124 -1459
rect 1390 -1528 1395 -1523
rect 120 -1541 125 -1536
rect 122 -1586 127 -1581
rect -19 -1615 -14 -1610
<< metal2 >>
rect 337 227 1470 231
rect 337 193 341 227
rect 648 36 652 227
rect 648 32 805 36
rect 89 -8 93 22
rect 648 1 652 32
rect -243 -12 93 -8
rect -243 -182 -239 -12
rect -4 -182 -1 -68
rect 113 -70 119 -31
rect 51 -76 119 -70
rect 51 -164 57 -76
rect 113 -112 119 -76
rect 442 -123 445 -81
rect 442 -126 606 -123
rect 442 -166 445 -126
rect 163 -167 445 -166
rect 158 -169 445 -167
rect -243 -186 -55 -182
rect -4 -185 216 -182
rect -243 -427 -239 -186
rect -59 -205 -55 -186
rect 257 -205 261 -169
rect -59 -209 261 -205
rect 442 -205 445 -169
rect 442 -208 533 -205
rect 54 -266 58 -228
rect 530 -320 533 -208
rect 624 -299 627 -85
rect 645 -307 649 -86
rect 663 -141 666 -86
rect 801 -100 805 32
rect 975 -34 1227 -31
rect 774 -122 922 -119
rect 774 -141 777 -122
rect 663 -144 777 -141
rect 724 -281 727 -246
rect 743 -307 747 -246
rect 761 -298 764 -247
rect 919 -298 922 -122
rect 1224 -159 1227 -34
rect 1466 -52 1470 227
rect 1391 -58 1591 -52
rect 1391 -112 1397 -58
rect 1224 -162 1342 -159
rect 1167 -170 1320 -167
rect 943 -194 960 -191
rect 761 -301 925 -298
rect 645 -311 747 -307
rect 530 -323 699 -320
rect 743 -394 747 -311
rect 743 -398 874 -394
rect 78 -427 82 -403
rect -243 -431 82 -427
rect -243 -1775 -239 -431
rect 487 -440 543 -436
rect 150 -445 306 -444
rect 487 -445 491 -440
rect 150 -448 491 -445
rect 150 -459 154 -448
rect 302 -449 491 -448
rect 539 -444 543 -440
rect 13 -645 16 -501
rect 109 -512 151 -509
rect 109 -546 112 -512
rect 109 -549 289 -546
rect 109 -604 112 -549
rect 302 -558 306 -449
rect 146 -561 481 -558
rect 146 -562 493 -561
rect 477 -565 493 -562
rect 13 -648 458 -645
rect -22 -668 146 -664
rect -22 -891 -18 -668
rect 477 -685 481 -565
rect 399 -689 481 -685
rect 512 -715 516 -501
rect 531 -538 534 -501
rect 531 -541 830 -538
rect 653 -715 657 -629
rect 672 -694 675 -628
rect 827 -694 830 -541
rect 870 -679 874 -398
rect 885 -466 901 -463
rect 922 -664 925 -301
rect 957 -496 960 -194
rect 1167 -463 1170 -170
rect 1317 -175 1320 -170
rect 1339 -175 1342 -162
rect 1298 -184 1301 -179
rect 1280 -187 1301 -184
rect 1280 -233 1283 -187
rect 1280 -236 1308 -233
rect 1305 -335 1308 -236
rect 1305 -338 1521 -335
rect 1000 -466 1170 -463
rect 1195 -448 1462 -445
rect 1195 -496 1198 -448
rect 957 -499 1198 -496
rect 1268 -586 1272 -549
rect 1289 -580 1292 -549
rect 1156 -590 1272 -586
rect 1156 -679 1160 -590
rect 1211 -612 1380 -609
rect 870 -683 1160 -679
rect 672 -697 1070 -694
rect 512 -719 657 -715
rect 401 -741 480 -737
rect 98 -891 102 -861
rect -22 -895 102 -891
rect 40 -1091 43 -965
rect 98 -976 102 -895
rect 476 -908 480 -741
rect 653 -751 657 -719
rect 653 -755 765 -751
rect 761 -792 765 -755
rect 1156 -792 1160 -683
rect 729 -796 1160 -792
rect 1377 -801 1380 -612
rect 1297 -804 1380 -801
rect 1297 -904 1300 -804
rect 1459 -853 1462 -448
rect 1345 -856 1462 -853
rect 1345 -905 1348 -856
rect 767 -932 773 -924
rect 767 -938 777 -932
rect 593 -955 596 -949
rect 593 -958 601 -955
rect 141 -976 145 -970
rect 84 -980 542 -976
rect 84 -1058 88 -980
rect 538 -990 542 -980
rect 538 -994 563 -990
rect 598 -996 601 -958
rect 771 -966 777 -938
rect 1518 -944 1521 -338
rect 1585 -463 1591 -58
rect 1646 -232 1702 -229
rect 1559 -469 1605 -463
rect 1183 -947 1521 -944
rect 771 -972 918 -966
rect 1599 -970 1605 -469
rect 1699 -569 1702 -232
rect 1665 -572 1704 -569
rect 771 -996 777 -972
rect 598 -999 618 -996
rect 40 -1094 540 -1091
rect 315 -1130 494 -1126
rect 315 -1150 319 -1130
rect 490 -1220 494 -1130
rect 615 -1168 618 -999
rect 912 -999 918 -972
rect 1401 -976 1605 -970
rect 1401 -999 1407 -976
rect 912 -1005 1407 -999
rect 1493 -1003 1499 -976
rect 764 -1168 767 -1077
rect 615 -1171 771 -1168
rect 615 -1185 618 -1171
rect 912 -1220 918 -1005
rect 1200 -1074 1392 -1071
rect 490 -1226 918 -1220
rect 1508 -1143 1511 -1117
rect 1508 -1146 1529 -1143
rect -35 -1612 -32 -1356
rect 65 -1504 68 -1322
rect 490 -1386 494 -1226
rect 266 -1390 494 -1386
rect 119 -1414 172 -1411
rect 124 -1416 172 -1414
rect 167 -1419 172 -1416
rect 167 -1424 244 -1419
rect 266 -1421 270 -1390
rect 319 -1442 374 -1437
rect 119 -1504 122 -1464
rect 65 -1507 122 -1504
rect 119 -1518 122 -1507
rect 247 -1518 250 -1502
rect 119 -1519 250 -1518
rect 96 -1521 250 -1519
rect 96 -1522 122 -1521
rect 96 -1589 99 -1522
rect 120 -1535 247 -1530
rect 120 -1536 125 -1535
rect 242 -1542 247 -1535
rect 369 -1538 374 -1442
rect 326 -1543 374 -1538
rect 122 -1589 125 -1586
rect 96 -1592 125 -1589
rect -35 -1615 -19 -1612
rect 111 -1639 114 -1592
rect 257 -1639 260 -1620
rect 111 -1642 260 -1639
rect 207 -1673 210 -1642
rect 553 -1673 556 -1245
rect 1390 -1523 1393 -1147
rect 1526 -1188 1529 -1146
rect 1701 -1188 1704 -572
rect 1526 -1191 1704 -1188
rect 1526 -1673 1529 -1191
rect 207 -1676 1529 -1673
rect 415 -1775 419 -1676
rect -243 -1779 419 -1775
use XNOR  XNOR_3
timestamp 1701464944
transform 1 0 -5 0 1 -1325
box -10 -18 447 179
use AND  AND_1
timestamp 1701359634
transform 1 0 242 0 1 -1618
box -2 -4 111 81
use AND  AND_0
timestamp 1701359634
transform 1 0 237 0 1 -1500
box -2 -4 111 81
use not  not_7
timestamp 1698047077
transform 1 0 129 0 1 -1561
box -9 -20 16 20
use not  not_6
timestamp 1698047077
transform 1 0 128 0 1 -1439
box -9 -20 16 20
use not  not_5
timestamp 1698047077
transform 1 0 149 0 1 -1042
box -9 -20 16 20
use not  not_4
timestamp 1698047077
transform 1 0 147 0 1 -945
box -9 -20 16 20
use AND3  AND3_1
timestamp 1701468290
transform 1 0 758 0 1 -1058
box -31 -53 128 22
use AND3  AND3_0
timestamp 1701468290
transform 1 0 588 0 1 -931
box -31 -53 128 22
use OR4  OR4_1
timestamp 1701474829
transform 1 0 1439 0 1 -1052
box -21 -61 154 41
use XNOR  XNOR_2
timestamp 1701464944
transform 1 0 -11 0 1 -864
box -10 -18 447 179
use not  not_3
timestamp 1698047077
transform 1 0 153 0 1 -587
box -9 -20 16 20
use AND4  AND4_2
timestamp 1701469746
transform 1 0 646 0 1 -612
box -27 -46 129 35
use AND4  AND4_0
timestamp 1701469746
transform 1 0 1257 0 1 -520
box -27 -46 129 35
use XNOR  XNOR_1
timestamp 1701464944
transform 1 0 1 0 1 -406
box -10 -18 447 179
use not  not_2
timestamp 1698047077
transform 1 0 153 0 1 -484
box -9 -20 16 20
use AND4  AND4_1
timestamp 1701469746
transform 1 0 504 0 1 -484
box -27 -46 129 35
use AND5  AND5_1
timestamp 1701473697
transform 1 0 710 0 1 -232
box -22 -45 148 78
use OR4  OR4_0
timestamp 1701474829
transform 1 0 1305 0 1 -157
box -21 -61 154 41
use XNOR  XNOR_0
timestamp 1701464944
transform 1 0 10 0 1 18
box -10 -18 447 179
use not  not_0
timestamp 1698047077
transform 1 0 151 0 1 -41
box -9 -20 16 20
use not  not_1
timestamp 1698047077
transform 1 0 153 0 1 -142
box -9 -20 16 20
use AND5  AND5_0
timestamp 1701473697
transform 1 0 612 0 1 -72
box -22 -45 148 78
<< labels >>
rlabel metal1 1409 -531 1412 -530 1 equal
rlabel metal1 1616 -1073 1619 -1072 1 lesser
rlabel metal1 -120 131 -117 132 1 A0
rlabel metal1 -79 42 -76 43 1 B0
rlabel metal1 -151 -293 -148 -292 1 A1
rlabel metal1 -59 -382 -56 -381 1 B1
rlabel metal1 -158 -750 -155 -749 1 A2
rlabel metal1 -74 -840 -71 -839 1 B2
rlabel metal1 -202 -1211 -199 -1210 1 A3
rlabel metal1 -95 -1301 -92 -1300 1 B3
rlabel metal2 426 228 431 229 5 vdd
rlabel metal2 181 -1778 186 -1777 1 gnd
rlabel metal1 1530 -178 1532 -177 1 greater
<< end >>
