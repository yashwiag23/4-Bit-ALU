magic
tech scmos
timestamp 1701365046
<< metal1 >>
rect 1044 465 1147 469
rect 5 202 78 209
rect 165 187 199 197
rect 1271 169 1373 172
rect -29 119 10 129
rect 1370 -321 1373 169
rect -226 -324 1373 -321
rect -226 -900 -223 -324
rect 1043 -900 1077 -896
rect -226 -1185 -222 -900
rect -37 -1163 78 -1156
rect 66 -1177 129 -1173
rect 66 -1185 70 -1177
rect 179 -1176 196 -1169
rect 179 -1177 187 -1176
rect -226 -1189 70 -1185
rect 1270 -1196 1345 -1193
rect -101 -1246 8 -1236
rect 1342 -1758 1345 -1196
rect -171 -1761 1345 -1758
rect -171 -2484 -168 -1761
rect 1027 -2210 1068 -2206
rect -25 -2473 63 -2466
rect -171 -2487 113 -2484
rect 155 -2486 179 -2480
rect 1252 -2506 1337 -2503
rect -73 -2556 -8 -2546
rect 1334 -3054 1337 -2506
rect -187 -3057 1337 -3054
rect -187 -3735 -184 -3057
rect 1043 -3440 1074 -3436
rect 11 -3703 78 -3696
rect 83 -3715 129 -3712
rect 173 -3715 195 -3710
rect 83 -3735 86 -3715
rect -187 -3738 86 -3735
rect 1271 -3736 1289 -3733
rect -35 -3786 8 -3776
<< m2contact >>
rect 129 -1179 135 -1173
rect 172 -1177 179 -1170
rect 113 -2487 118 -2482
rect 149 -2486 155 -2480
rect 129 -3715 134 -3710
rect 168 -3715 173 -3710
<< metal2 >>
rect 472 693 1643 698
rect 472 561 477 693
rect 464 -213 472 6
rect -406 -221 472 -213
rect -406 -1635 -398 -221
rect 1638 -563 1643 693
rect 481 -568 1643 -563
rect 481 -802 486 -568
rect 135 -1177 172 -1173
rect 409 -1635 417 -1357
rect -406 -1643 417 -1635
rect -406 -2897 -398 -1643
rect 1638 -1878 1643 -568
rect 490 -1883 1643 -1878
rect 490 -2113 495 -1883
rect 145 -2482 149 -2481
rect 118 -2486 149 -2482
rect 443 -2897 451 -2671
rect -406 -2905 451 -2897
rect -406 -4133 -398 -2905
rect 1638 -3187 1643 -1883
rect 447 -3192 1643 -3187
rect 447 -3342 452 -3192
rect 134 -3715 168 -3710
rect 412 -4133 420 -3897
rect -406 -4141 420 -4133
use fulladder  fulladder_0
timestamp 1701362989
transform 1 0 167 0 1 284
box -167 -284 1109 282
use fulladder  fulladder_1
timestamp 1701362989
transform 1 0 165 0 1 -1081
box -167 -284 1109 282
use fulladder  fulladder_2
timestamp 1701362989
transform 1 0 149 0 1 -2391
box -167 -284 1109 282
use fulladder  fulladder_3
timestamp 1701362989
transform 1 0 165 0 1 -3621
box -167 -284 1109 282
<< labels >>
rlabel metal1 167 188 172 193 1 Cin
rlabel metal1 -26 121 -24 126 1 B0
rlabel metal1 7 203 11 207 1 A0
rlabel metal2 849 694 856 697 5 vdd
rlabel metal2 123 -4139 134 -4135 1 gnd
rlabel metal1 1144 466 1146 467 1 S0
rlabel metal1 1074 -899 1076 -898 1 S1
rlabel metal1 1071 -3439 1073 -3437 1 S3
rlabel metal1 1287 -3735 1288 -3734 1 Cout
rlabel metal1 -35 -1161 -29 -1159 1 A1
rlabel metal1 -97 -1239 -91 -1237 1 B1
rlabel metal1 -24 -2471 -18 -2467 1 A2
rlabel metal1 -69 -2552 -65 -2549 1 B2
rlabel metal1 13 -3701 17 -3698 1 A3
rlabel metal1 -33 -3783 -28 -3779 1 B3
rlabel metal1 1062 -2209 1067 -2208 1 S2
<< end >>
