magic
tech scmos
timestamp 1701538289
<< metal1 >>
rect -89 66 -59 72
rect -62 30 -59 66
rect -62 27 3 30
rect -62 -88 -59 27
rect 18 22 21 30
rect 110 23 124 26
rect -23 19 21 22
rect -62 -91 4 -88
rect -62 -225 -59 -91
rect 19 -95 22 -88
rect 110 -95 122 -92
rect -15 -98 22 -95
rect -62 -228 4 -225
rect -62 -355 -59 -228
rect 19 -232 22 -225
rect 109 -232 130 -229
rect -14 -235 22 -232
rect -62 -358 4 -355
rect -62 -483 -59 -358
rect 19 -363 22 -355
rect 109 -362 131 -359
rect -9 -366 22 -363
rect -62 -486 6 -483
rect -62 -603 -59 -486
rect 20 -489 23 -483
rect -16 -492 23 -489
rect 108 -490 129 -487
rect -62 -606 7 -603
rect -62 -734 -59 -606
rect 22 -611 25 -603
rect 113 -610 139 -607
rect -20 -614 25 -611
rect -62 -737 5 -734
rect -62 -854 -59 -737
rect 20 -742 23 -734
rect 111 -741 141 -738
rect -23 -745 23 -742
rect -62 -857 3 -854
rect 21 -861 24 -854
rect 111 -861 153 -858
rect -22 -864 24 -861
<< metal2 >>
rect 84 115 175 120
rect 84 80 89 115
rect 16 -8 21 2
rect -32 -13 21 -8
rect -30 -124 -25 -13
rect 170 -33 175 115
rect 79 -38 175 -33
rect 19 -124 24 -113
rect -30 -129 24 -124
rect -30 -270 -25 -129
rect 170 -170 175 -38
rect 73 -175 175 -170
rect 15 -270 20 -250
rect -31 -275 20 -270
rect -30 -403 -25 -275
rect 170 -300 175 -175
rect 77 -305 175 -300
rect 16 -403 21 -380
rect -30 -408 21 -403
rect -30 -528 -25 -408
rect 170 -428 175 -305
rect 83 -433 175 -428
rect 19 -528 24 -508
rect -30 -533 24 -528
rect -30 -643 -25 -533
rect 170 -548 175 -433
rect 84 -553 175 -548
rect -29 -646 -25 -643
rect 32 -646 37 -628
rect -29 -651 37 -646
rect -29 -657 -25 -651
rect -30 -782 -25 -657
rect 170 -679 175 -553
rect 85 -684 175 -679
rect 16 -782 21 -759
rect -30 -787 21 -782
rect -30 -911 -25 -787
rect 170 -799 175 -684
rect 85 -804 175 -799
rect 13 -911 18 -879
rect -31 -916 18 -911
use AND  AND_0
timestamp 1701359634
transform 1 0 2 0 1 4
box -2 -4 111 81
use AND  AND_1
timestamp 1701359634
transform 1 0 3 0 1 -114
box -2 -4 111 81
use AND  AND_2
timestamp 1701359634
transform 1 0 3 0 1 -251
box -2 -4 111 81
use AND  AND_3
timestamp 1701359634
transform 1 0 3 0 1 -381
box -2 -4 111 81
use AND  AND_4
timestamp 1701359634
transform 1 0 4 0 1 -509
box -2 -4 111 81
use AND  AND_5
timestamp 1701359634
transform 1 0 6 0 1 -629
box -2 -4 111 81
use AND  AND_6
timestamp 1701359634
transform 1 0 4 0 1 -760
box -2 -4 111 81
use AND  AND_7
timestamp 1701359634
transform 1 0 5 0 1 -880
box -2 -4 111 81
<< labels >>
rlabel metal2 117 116 121 118 5 vdd
rlabel space -33 -914 -28 -913 1 gnd
rlabel metal1 -82 68 -78 70 1 enable
rlabel metal1 -20 20 -16 22 1 A0
rlabel metal1 -12 -97 -8 -95 1 A1
rlabel metal1 -11 -234 -10 -233 1 A2
rlabel metal1 -7 -365 -6 -364 1 A3
rlabel metal1 -12 -491 -11 -490 1 B0
rlabel metal1 -16 -613 -15 -612 1 B1
rlabel metal1 -18 -744 -17 -743 1 B2
rlabel metal1 -18 -863 -17 -862 1 B3
rlabel metal1 120 24 122 25 1 F0
rlabel metal1 119 -94 121 -93 1 F1
rlabel metal1 126 -231 128 -230 1 F2
rlabel metal1 127 -361 129 -360 1 F3
rlabel metal1 125 -489 127 -488 1 F4
rlabel metal1 134 -609 136 -608 1 F5
rlabel metal1 137 -740 139 -739 1 F6
rlabel metal1 147 -860 149 -859 1 F7
<< end >>
