magic
tech scmos
timestamp 1701474829
<< nwell >>
rect -21 0 66 21
<< ntransistor >>
rect -10 -45 -8 -39
rect 8 -45 10 -39
rect 28 -45 30 -39
rect 48 -45 50 -39
<< ptransistor >>
rect -10 9 -8 14
rect 8 9 10 14
rect 28 9 30 14
rect 48 9 50 14
<< ndiffusion >>
rect -12 -45 -10 -39
rect -8 -45 -7 -39
rect 5 -45 8 -39
rect 10 -45 12 -39
rect 24 -45 28 -39
rect 30 -45 33 -39
rect 45 -45 48 -39
rect 50 -45 53 -39
<< pdiffusion >>
rect -11 9 -10 14
rect -8 9 8 14
rect 10 9 28 14
rect 30 9 48 14
rect 50 9 52 14
<< ndcontact >>
rect -16 -45 -12 -39
rect -7 -45 -3 -39
rect 1 -45 5 -39
rect 12 -45 16 -39
rect 20 -45 24 -39
rect 33 -45 37 -39
rect 41 -45 45 -39
rect 53 -45 57 -39
<< pdcontact >>
rect -15 9 -11 14
rect 52 9 56 14
<< polysilicon >>
rect -10 14 -8 17
rect 8 14 10 17
rect 28 14 30 17
rect 48 14 50 18
rect -10 -17 -8 9
rect 8 -17 10 9
rect -13 -21 -8 -17
rect 5 -21 10 -17
rect 28 -19 30 9
rect 48 -18 50 9
rect -10 -39 -8 -21
rect 8 -39 10 -21
rect 24 -23 30 -19
rect 46 -22 50 -18
rect 28 -39 30 -23
rect 48 -39 50 -22
rect -10 -50 -8 -45
rect 8 -50 10 -45
rect 28 -50 30 -45
rect 48 -50 50 -45
<< polycontact >>
rect -17 -21 -13 -17
rect 1 -21 5 -17
rect 20 -23 24 -19
rect 42 -22 46 -18
<< metal1 >>
rect 36 40 42 41
rect 36 37 126 40
rect 36 27 42 37
rect -21 21 66 27
rect -15 14 -12 21
rect -21 -21 -17 -17
rect -3 -21 1 -17
rect 16 -23 20 -19
rect 38 -22 42 -18
rect 53 -21 56 9
rect 123 2 126 37
rect 104 -21 118 -19
rect 53 -22 118 -21
rect 138 -22 154 -19
rect 53 -24 107 -22
rect 53 -33 56 -24
rect -6 -36 56 -33
rect -6 -39 -3 -36
rect 13 -39 16 -36
rect 34 -39 37 -36
rect 53 -39 56 -36
rect -16 -57 -12 -45
rect 2 -50 5 -45
rect 0 -53 5 -50
rect 0 -57 3 -53
rect 20 -57 23 -45
rect 41 -57 44 -45
rect 118 -48 121 -35
rect 102 -51 121 -48
rect 102 -57 105 -51
rect -16 -60 105 -57
rect -16 -61 -12 -60
use not  not_0
timestamp 1698047077
transform 1 0 125 0 1 -17
box -9 -20 16 20
<< labels >>
rlabel metal1 151 -21 152 -20 7 out
rlabel metal1 82 -59 83 -58 1 gnd
rlabel metal1 40 -20 41 -19 1 D
rlabel metal1 17 -21 18 -20 1 C
rlabel metal1 -2 -20 -1 -19 1 B
rlabel metal1 -20 -20 -19 -19 3 A
rlabel metal1 38 32 39 33 1 vdd
<< end >>
