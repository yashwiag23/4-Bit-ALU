* NGSPICE file created from decoder.ext - technology: scmos

.global Vdd Gnd 

.subckt NAND gnd A B out vdd
M1000 a_13_n30# A gnd Gnd nfet w=3u l=1.2u
+  ad=28.8p pd=25.2u as=21.6p ps=20.4u
M1001 out B a_13_n30# Gnd nfet w=3u l=1.2u
+  ad=14.4p pd=15.6u as=0p ps=0u
M1002 out B vdd w_n1_n1# pfet w=2.4u l=1.2u
+  ad=14.4p pd=21.6u as=17.28p ps=24u
M1003 out A vdd w_n1_n1# pfet w=2.4u l=1.2u
+  ad=0p pd=0u as=0p ps=0u
.ends

.subckt not gnd VDD in out
M1000 out in gnd Gnd nfet w=2.4u l=1.2u
+  ad=7.2p pd=10.8u as=7.2p ps=10.8u
M1001 out in VDD w_n9_1# pfet w=2.4u l=1.2u
+  ad=7.2p pd=10.8u as=7.2p ps=10.8u
.ends

.subckt AND gnd A B out vdd
XNAND_0 gnd A B not_0/in vdd NAND
Xnot_0 gnd vdd not_0/in out not
.ends


* Top level circuit decoder

XAND_1 gnd s0 AND_1/B en1 vdd AND
XAND_0 gnd AND_2/B AND_1/B en0 vdd AND
XAND_2 gnd s1 AND_2/B en2 vdd AND
Xnot_0 gnd vdd s0 AND_2/B not
XAND_3 gnd s1 s0 en3 vdd AND
Xnot_1 gnd vdd s1 AND_1/B not
.end

